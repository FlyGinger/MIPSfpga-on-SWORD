// Author: Jiang Zengkai
// Date: 2019.5.18

module io_sd(
    input wire clk, // 100 MHz
    input wire rst, // reset, active high
    output wire sd_clk,
    input wire sd_cd, // card detect, not used
    inout wire sd_cmd, // command
    inout wire [3:0] sd_dat // data
);

    // SD card clock generation
    






endmodule