// Author: Jiang Zengkai
// Date: 2019.3.21
// Version: 1.0

module clk_div(
    input wire clk, // 50 MHz
    output reg [31:0] clk_div);
    
    always @ (posedge clk) begin
        clk_div <= clk_div + 1;
    end

endmodule

// 0: 25 MHz
// 1: 12.5 MHz
// 2: 6.25 MHz
// 3: 3.125 MHz
// 4: 1.5625 MHz
// 5: 781.25 KHz
// 6: 390.625 KHz
// 7: 195.53125 KHz
// 8: 97.65625 KHz
// 9: 48.828125 KHz
// 10: 24.4140625 KHz
// 11: 12.2070313 KHz
// 12: 6.10351565 KHz
// 13: 3.05175783 KHz
// 14: 1.52587892 KHz
// 15: 762.93946 Hz
// 16: 381.46973 Hz
// 17: 190.734865 Hz
// 18: 95.3674325 Hz
// 19: 47.6837163 Hz
// 20: 23.8418582 Hz
// 21: 11.9209291 Hz
// 22: 5.96046455 Hz
// 23: 2.98023228 Hz
// 24: 1.49011614 Hz
// 25: 1/(1.34s)
// 26: 1/(2.68s)
// 27: 1/(5.37s)
// 28: 1/(10.74s)
// 29: 1/(21.47s)
// 30: 1/(42.95s)
// 31: 1/(85.90s)
